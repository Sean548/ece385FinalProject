//create collision detection and what happens based on the type of the objects when they collide